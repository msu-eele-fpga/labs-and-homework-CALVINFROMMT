library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.std_logic_unsigned.all;


entity hps_led_control is
	port();

end entity;

architecture hps_led_control_arch of hps_led_control is 

begin



end architecture;